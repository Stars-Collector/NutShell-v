//commit 5dafedae3450c366c2197a53bbdce14726fbe194
//Merge: d114ea0 ecce4b9
//Author: Yinan Xu <xuyinan@ict.ac.cn>
//Date:   Mon Aug 26 09:50:32 2024 +0800
//
//    Merge pull request #206 from zhangziqing/oscpu-master-wip
//    
//    NutShell master branch re-adaption for FPGA platforms
//diff --git a/Makefile b/Makefile
//index ad28764..c34d99d 100644
//--- a/Makefile
//+++ b/Makefile
//@@ -19,7 +19,7 @@ SIMTOP = top.TopMain
// IMAGE ?= ready-to-run/linux.bin
// 
// DATAWIDTH ?= 64
//-BOARD ?= sim  # sim  pynq  axu3cg
//+BOARD ?= pynq  # sim  pynq  axu3cg
// CORE  ?= inorder  # inorder  ooo  embedded
// 
// MILL_ARGS_ALL  = $(MILL_ARGS)
//diff --git a/debian_on_fpga.gif b/debian_on_fpga.gif
//deleted file mode 100755
//index 8ae9ec2..0000000
//Binary files a/debian_on_fpga.gif and /dev/null differ
// Generated by CIRCT firtool-1.62.0
// Standard header to adapt well known macros for register randomization.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for prints and assertions.

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module Top(	// src/test/scala/TopMain.scala:28:7
  input clock,	// src/test/scala/TopMain.scala:28:7
        reset	// src/test/scala/TopMain.scala:28:7
);

  NutShell nutshell (	// src/test/scala/TopMain.scala:30:24
    .clock                     (clock),
    .reset                     (reset),
    .io_mem_awready           (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_awvalid           (/* unused */),
    .io_mem_awaddr       (/* unused */),
    .io_mem_awprot       (/* unused */),
    .io_mem_awid         (/* unused */),
    .io_mem_awuser       (/* unused */),
    .io_mem_awlen        (/* unused */),
    .io_mem_awsize       (/* unused */),
    .io_mem_awburst      (/* unused */),
    .io_mem_awlock       (/* unused */),
    .io_mem_awcache      (/* unused */),
    .io_mem_awqos        (/* unused */),
    .io_mem_wready            (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_wvalid            (/* unused */),
    .io_mem_wdata        (/* unused */),
    .io_mem_wstrb        (/* unused */),
    .io_mem_wlast        (/* unused */),
    .io_mem_bready            (/* unused */),
    .io_mem_bvalid            (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_bresp        (2'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_bid          (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_buser        (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_arready           (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_arvalid           (/* unused */),
    .io_mem_araddr       (/* unused */),
    .io_mem_arprot       (/* unused */),
    .io_mem_arid         (/* unused */),
    .io_mem_aruser       (/* unused */),
    .io_mem_arlen        (/* unused */),
    .io_mem_arsize       (/* unused */),
    .io_mem_arburst      (/* unused */),
    .io_mem_arlock       (/* unused */),
    .io_mem_arcache      (/* unused */),
    .io_mem_arqos        (/* unused */),
    .io_mem_rready            (/* unused */),
    .io_mem_rvalid            (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_rresp        (2'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_rdata        (64'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_rlast        (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_rid          (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mem_ruser        (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_awready          (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_awvalid          (/* unused */),
    .io_mmio_awaddr      (/* unused */),
    .io_mmio_awprot      (/* unused */),
    .io_mmio_awid        (/* unused */),
    .io_mmio_awuser      (/* unused */),
    .io_mmio_awlen       (/* unused */),
    .io_mmio_awsize      (/* unused */),
    .io_mmio_awburst     (/* unused */),
    .io_mmio_awlock      (/* unused */),
    .io_mmio_awcache     (/* unused */),
    .io_mmio_awqos       (/* unused */),
    .io_mmio_wready           (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_wvalid           (/* unused */),
    .io_mmio_wdata       (/* unused */),
    .io_mmio_wstrb       (/* unused */),
    .io_mmio_wlast       (/* unused */),
    .io_mmio_bready           (/* unused */),
    .io_mmio_bvalid           (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_bresp       (2'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_bid         (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_buser       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_arready          (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_arvalid          (/* unused */),
    .io_mmio_araddr      (/* unused */),
    .io_mmio_arprot      (/* unused */),
    .io_mmio_arid        (/* unused */),
    .io_mmio_aruser      (/* unused */),
    .io_mmio_arlen       (/* unused */),
    .io_mmio_arsize      (/* unused */),
    .io_mmio_arburst     (/* unused */),
    .io_mmio_arlock      (/* unused */),
    .io_mmio_arcache     (/* unused */),
    .io_mmio_arqos       (/* unused */),
    .io_mmio_rready           (/* unused */),
    .io_mmio_rvalid           (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_rresp       (2'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_rdata       (64'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_rlast       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_rid         (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_mmio_ruser       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awready      (/* unused */),
    .io_frontend_awvalid      (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awaddr  (32'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awprot  (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awid    (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awuser  (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awlen   (8'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awsize  (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awburst (2'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awlock  (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awcache (4'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_awqos   (4'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_wready       (/* unused */),
    .io_frontend_wvalid       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_wdata   (64'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_wstrb   (8'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_wlast   (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_bready       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_bvalid       (/* unused */),
    .io_frontend_bresp   (/* unused */),
    .io_frontend_bid     (/* unused */),
    .io_frontend_buser   (/* unused */),
    .io_frontend_arready      (/* unused */),
    .io_frontend_arvalid      (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_araddr  (32'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arprot  (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arid    (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_aruser  (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arlen   (8'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arsize  (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arburst (2'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arlock  (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arcache (4'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_arqos   (4'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_rready       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_frontend_rvalid       (/* unused */),
    .io_frontend_rresp   (/* unused */),
    .io_frontend_rdata   (/* unused */),
    .io_frontend_rlast   (/* unused */),
    .io_frontend_rid     (/* unused */),
    .io_frontend_ruser   (/* unused */),
    .io_meip                   (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_ila_WBUpc              (/* unused */),
    .io_ila_WBUvalid           (/* unused */),
    .io_ila_WBUrfWen           (/* unused */),
    .io_ila_WBUrfDest          (/* unused */),
    .io_ila_WBUrfData          (/* unused */),
    .io_ila_InstrCnt           (/* unused */)
  );
  AXI4VGA vga (	// src/test/scala/TopMain.scala:31:19
    .clock                   (clock),
    .reset                   (reset),
    .io_in_fb_awready       (/* unused */),
    .io_in_fb_awvalid       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_awaddr   (32'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_awprot   (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_wready        (/* unused */),
    .io_in_fb_wvalid        (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_wdata    (64'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_wstrb    (8'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_bready        (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_bvalid        (/* unused */),
    .io_in_fb_bresp    (/* unused */),
    .io_in_fb_arready       (/* unused */),
    .io_in_fb_arvalid       (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_araddr   (32'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_arprot   (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_rready        (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_fb_rvalid        (/* unused */),
    .io_in_fb_rresp    (/* unused */),
    .io_in_fb_rdata    (/* unused */),
    .io_in_ctrl_awready     (/* unused */),
    .io_in_ctrl_awvalid     (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_awaddr (32'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_awprot (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_wready      (/* unused */),
    .io_in_ctrl_wvalid      (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_wdata  (64'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_wstrb  (8'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_bready      (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_bvalid      (/* unused */),
    .io_in_ctrl_bresp  (/* unused */),
    .io_in_ctrl_arready     (/* unused */),
    .io_in_ctrl_arvalid     (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_araddr (32'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_arprot (3'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_rready      (1'h0),	// src/test/scala/TopMain.scala:33:15
    .io_in_ctrl_rvalid      (/* unused */),
    .io_in_ctrl_rresp  (/* unused */),
    .io_in_ctrl_rdata  (/* unused */),
    .io_vga_rgb              (/* unused */),
    .io_vga_hsync            (/* unused */),
    .io_vga_vsync            (/* unused */),
    .io_vga_valid            (/* unused */)
  );
endmodule

