//commit 5dafedae3450c366c2197a53bbdce14726fbe194
//Merge: d114ea0 ecce4b9
//Author: Yinan Xu <xuyinan@ict.ac.cn>
//Date:   Mon Aug 26 09:50:32 2024 +0800
//
//    Merge pull request #206 from zhangziqing/oscpu-master-wip
//    
//    NutShell master branch re-adaption for FPGA platforms
//diff --git a/debian_on_fpga.gif b/debian_on_fpga.gif
//deleted file mode 100755
//index 8ae9ec2..0000000
//Binary files a/debian_on_fpga.gif and /dev/null differ
// Generated by CIRCT firtool-1.62.0
// Standard header to adapt well known macros for register randomization.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for prints and assertions.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module SimTop(	// src/main/scala/sim/NutShellSim.scala:26:7
  input         clock,	// src/main/scala/sim/NutShellSim.scala:26:7
                reset,	// src/main/scala/sim/NutShellSim.scala:26:7
  output [63:0] difftest_step,	// difftest/src/main/scala/Difftest.scala:393:22
  input         difftest_perfCtrl_clean,	// difftest/src/main/scala/Difftest.scala:393:22
                difftest_perfCtrl_dump,	// difftest/src/main/scala/Difftest.scala:393:22
  input  [63:0] difftest_logCtrl_begin,	// difftest/src/main/scala/Difftest.scala:393:22
                difftest_logCtrl_end,	// difftest/src/main/scala/Difftest.scala:393:22
                difftest_logCtrl_level,	// difftest/src/main/scala/Difftest.scala:393:22
  output        difftest_uart_out_valid,	// difftest/src/main/scala/Difftest.scala:393:22
  output [7:0]  difftest_uart_out_ch,	// difftest/src/main/scala/Difftest.scala:393:22
  output        difftest_uart_in_valid,	// difftest/src/main/scala/Difftest.scala:393:22
  input  [7:0]  difftest_uart_in_ch	// difftest/src/main/scala/Difftest.scala:393:22
);

  wire        _mmio_io_rw_req_ready;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_rw_resp_valid;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire [3:0]  _mmio_io_rw_resp_bits_cmd;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire [63:0] _mmio_io_rw_resp_bits_rdata;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_meip;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_dma_awvalid;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire [31:0] _mmio_io_dma_awaddr;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_dma_wvalid;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire [63:0] _mmio_io_dma_wdata;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire [7:0]  _mmio_io_dma_wstrb;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_dma_bready;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_dma_arvalid;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire [31:0] _mmio_io_dma_araddr;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _mmio_io_dma_rready;	// src/main/scala/sim/NutShellSim.scala:33:20
  wire        _memdelay_io_in_awready;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_in_wready;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_in_bvalid;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_in_arready;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_in_rvalid;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire [63:0] _memdelay_io_in_rdata;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_in_rlast;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_out_awvalid;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire [31:0] _memdelay_io_out_awaddr;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_out_wvalid;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire [63:0] _memdelay_io_out_wdata;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_out_wlast;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _memdelay_io_out_arvalid;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire [31:0] _memdelay_io_out_araddr;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire [7:0]  _memdelay_io_out_arlen;	// src/main/scala/sim/NutShellSim.scala:32:24
  wire        _mem_io_in_awready;	// src/main/scala/sim/NutShellSim.scala:29:19
  wire        _mem_io_in_wready;	// src/main/scala/sim/NutShellSim.scala:29:19
  wire        _mem_io_in_bvalid;	// src/main/scala/sim/NutShellSim.scala:29:19
  wire        _mem_io_in_rvalid;	// src/main/scala/sim/NutShellSim.scala:29:19
  wire [63:0] _mem_io_in_rdata;	// src/main/scala/sim/NutShellSim.scala:29:19
  wire        _mem_io_in_rlast;	// src/main/scala/sim/NutShellSim.scala:29:19
  wire        _soc_io_mem_awvalid;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [31:0] _soc_io_mem_awaddr;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [7:0]  _soc_io_mem_awlen;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_mem_wvalid;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [63:0] _soc_io_mem_wdata;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_mem_wlast;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_mem_arvalid;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [31:0] _soc_io_mem_araddr;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [7:0]  _soc_io_mem_arlen;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_mmio_req_valid;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [31:0] _soc_io_mmio_req_bits_addr;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [2:0]  _soc_io_mmio_req_bits_size;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [3:0]  _soc_io_mmio_req_bits_cmd;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [7:0]  _soc_io_mmio_req_bits_wmask;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [63:0] _soc_io_mmio_req_bits_wdata;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_mmio_resp_ready;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_frontend_awready;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_frontend_wready;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_frontend_bvalid;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_frontend_arready;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire        _soc_io_frontend_rvalid;	// src/main/scala/sim/NutShellSim.scala:28:19
  wire [63:0] _soc_io_frontend_rdata;	// src/main/scala/sim/NutShellSim.scala:28:19
  reg  [63:0] difftest_timer;	// difftest/src/main/scala/Difftest.scala:397:24
  wire        difftest_log_enable =
    difftest_timer >= difftest_logCtrl_begin & difftest_timer < difftest_logCtrl_end;	// difftest/src/main/scala/Difftest.scala:397:24, :570:22, :571:{17,26,35}
  always @(posedge clock) begin	// src/main/scala/sim/NutShellSim.scala:26:7
    if (reset)	// src/main/scala/sim/NutShellSim.scala:26:7
      difftest_timer <= 64'h0;	// difftest/src/main/scala/Difftest.scala:397:24
    else	// src/main/scala/sim/NutShellSim.scala:26:7
      difftest_timer <= difftest_timer + 64'h1;	// difftest/src/main/scala/Difftest.scala:395:19, :397:24, :398:20
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_	// src/main/scala/sim/NutShellSim.scala:26:7
    `ifdef FIRRTL_BEFORE_INITIAL	// src/main/scala/sim/NutShellSim.scala:26:7
      `FIRRTL_BEFORE_INITIAL	// src/main/scala/sim/NutShellSim.scala:26:7
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin	// src/main/scala/sim/NutShellSim.scala:26:7
      automatic logic [31:0] _RANDOM[0:1];	// src/main/scala/sim/NutShellSim.scala:26:7
      `ifdef INIT_RANDOM_PROLOG_	// src/main/scala/sim/NutShellSim.scala:26:7
        `INIT_RANDOM_PROLOG_	// src/main/scala/sim/NutShellSim.scala:26:7
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT	// src/main/scala/sim/NutShellSim.scala:26:7
        for (logic [1:0] i = 2'h0; i < 2'h2; i += 2'h1) begin
          _RANDOM[i[0]] = `RANDOM;	// src/main/scala/sim/NutShellSim.scala:26:7
        end	// src/main/scala/sim/NutShellSim.scala:26:7
        difftest_timer = {_RANDOM[1'h0], _RANDOM[1'h1]};	// difftest/src/main/scala/Difftest.scala:397:24, src/main/scala/sim/NutShellSim.scala:26:7
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL	// src/main/scala/sim/NutShellSim.scala:26:7
      `FIRRTL_AFTER_INITIAL	// src/main/scala/sim/NutShellSim.scala:26:7
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  NutShell soc (	// src/main/scala/sim/NutShellSim.scala:28:19
    .clock                    (clock),
    .reset                    (reset),
    .io_mem_awready          (_memdelay_io_in_awready),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mem_awvalid          (_soc_io_mem_awvalid),
    .io_mem_awaddr      (_soc_io_mem_awaddr),
    .io_mem_awlen       (_soc_io_mem_awlen),
    .io_mem_wready           (_memdelay_io_in_wready),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mem_wvalid           (_soc_io_mem_wvalid),
    .io_mem_wdata       (_soc_io_mem_wdata),
    .io_mem_wlast       (_soc_io_mem_wlast),
    .io_mem_bvalid           (_memdelay_io_in_bvalid),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mem_arready          (_memdelay_io_in_arready),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mem_arvalid          (_soc_io_mem_arvalid),
    .io_mem_araddr      (_soc_io_mem_araddr),
    .io_mem_arlen       (_soc_io_mem_arlen),
    .io_mem_rvalid           (_memdelay_io_in_rvalid),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mem_rdata       (_memdelay_io_in_rdata),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mem_rlast       (_memdelay_io_in_rlast),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_mmio_req_ready        (_mmio_io_rw_req_ready),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_mmio_req_valid        (_soc_io_mmio_req_valid),
    .io_mmio_req_bits_addr    (_soc_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size    (_soc_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd     (_soc_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask   (_soc_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata   (_soc_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready       (_soc_io_mmio_resp_ready),
    .io_mmio_resp_valid       (_mmio_io_rw_resp_valid),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_mmio_resp_bits_cmd    (_mmio_io_rw_resp_bits_cmd),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_mmio_resp_bits_rdata  (_mmio_io_rw_resp_bits_rdata),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_awready     (_soc_io_frontend_awready),
    .io_frontend_awvalid     (_mmio_io_dma_awvalid),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_awaddr (_mmio_io_dma_awaddr),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_wready      (_soc_io_frontend_wready),
    .io_frontend_wvalid      (_mmio_io_dma_wvalid),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_wdata  (_mmio_io_dma_wdata),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_wstrb  (_mmio_io_dma_wstrb),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_bready      (_mmio_io_dma_bready),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_bvalid      (_soc_io_frontend_bvalid),
    .io_frontend_arready     (_soc_io_frontend_arready),
    .io_frontend_arvalid     (_mmio_io_dma_arvalid),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_araddr (_mmio_io_dma_araddr),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_rready      (_mmio_io_dma_rready),	// src/main/scala/sim/NutShellSim.scala:33:20
    .io_frontend_rvalid      (_soc_io_frontend_rvalid),
    .io_frontend_rdata  (_soc_io_frontend_rdata),
    .io_meip                  (_mmio_io_meip)	// src/main/scala/sim/NutShellSim.scala:33:20
  );
  AXI4RAM mem (	// src/main/scala/sim/NutShellSim.scala:29:19
    .clock              (clock),
    .reset              (reset),
    .io_in_awready     (_mem_io_in_awready),
    .io_in_awvalid     (_memdelay_io_out_awvalid),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_awaddr (_memdelay_io_out_awaddr),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_wready      (_mem_io_in_wready),
    .io_in_wvalid      (_memdelay_io_out_wvalid),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_wdata  (_memdelay_io_out_wdata),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_wlast  (_memdelay_io_out_wlast),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_bvalid      (_mem_io_in_bvalid),
    .io_in_arvalid     (_memdelay_io_out_arvalid),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_araddr (_memdelay_io_out_araddr),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_arlen  (_memdelay_io_out_arlen),	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_rvalid      (_mem_io_in_rvalid),
    .io_in_rdata  (_mem_io_in_rdata),
    .io_in_rlast  (_mem_io_in_rlast)
  );
  AXI4Delayer memdelay (	// src/main/scala/sim/NutShellSim.scala:32:24
    .io_in_awready      (_memdelay_io_in_awready),
    .io_in_awvalid      (_soc_io_mem_awvalid),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_awaddr  (_soc_io_mem_awaddr),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_awlen   (_soc_io_mem_awlen),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_wready       (_memdelay_io_in_wready),
    .io_in_wvalid       (_soc_io_mem_wvalid),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_wdata   (_soc_io_mem_wdata),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_wlast   (_soc_io_mem_wlast),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_bvalid       (_memdelay_io_in_bvalid),
    .io_in_arready      (_memdelay_io_in_arready),
    .io_in_arvalid      (_soc_io_mem_arvalid),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_araddr  (_soc_io_mem_araddr),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_arlen   (_soc_io_mem_arlen),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_in_rvalid       (_memdelay_io_in_rvalid),
    .io_in_rdata   (_memdelay_io_in_rdata),
    .io_in_rlast   (_memdelay_io_in_rlast),
    .io_out_awready     (_mem_io_in_awready),	// src/main/scala/sim/NutShellSim.scala:29:19
    .io_out_awvalid     (_memdelay_io_out_awvalid),
    .io_out_awaddr (_memdelay_io_out_awaddr),
    .io_out_wready      (_mem_io_in_wready),	// src/main/scala/sim/NutShellSim.scala:29:19
    .io_out_wvalid      (_memdelay_io_out_wvalid),
    .io_out_wdata  (_memdelay_io_out_wdata),
    .io_out_wlast  (_memdelay_io_out_wlast),
    .io_out_bvalid      (_mem_io_in_bvalid),	// src/main/scala/sim/NutShellSim.scala:29:19
    .io_out_arvalid     (_memdelay_io_out_arvalid),
    .io_out_araddr (_memdelay_io_out_araddr),
    .io_out_arlen  (_memdelay_io_out_arlen),
    .io_out_rvalid      (_mem_io_in_rvalid),	// src/main/scala/sim/NutShellSim.scala:29:19
    .io_out_rdata  (_mem_io_in_rdata),	// src/main/scala/sim/NutShellSim.scala:29:19
    .io_out_rlast  (_mem_io_in_rlast)	// src/main/scala/sim/NutShellSim.scala:29:19
  );
  SimMMIO mmio (	// src/main/scala/sim/NutShellSim.scala:33:20
    .clock                 (clock),
    .reset                 (reset),
    .io_rw_req_ready       (_mmio_io_rw_req_ready),
    .io_rw_req_valid       (_soc_io_mmio_req_valid),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_req_bits_addr   (_soc_io_mmio_req_bits_addr),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_req_bits_size   (_soc_io_mmio_req_bits_size),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_req_bits_cmd    (_soc_io_mmio_req_bits_cmd),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_req_bits_wmask  (_soc_io_mmio_req_bits_wmask),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_req_bits_wdata  (_soc_io_mmio_req_bits_wdata),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_resp_ready      (_soc_io_mmio_resp_ready),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_rw_resp_valid      (_mmio_io_rw_resp_valid),
    .io_rw_resp_bits_cmd   (_mmio_io_rw_resp_bits_cmd),
    .io_rw_resp_bits_rdata (_mmio_io_rw_resp_bits_rdata),
    .io_meip               (_mmio_io_meip),
    .io_dma_awready       (_soc_io_frontend_awready),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_dma_awvalid       (_mmio_io_dma_awvalid),
    .io_dma_awaddr   (_mmio_io_dma_awaddr),
    .io_dma_wready        (_soc_io_frontend_wready),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_dma_wvalid        (_mmio_io_dma_wvalid),
    .io_dma_wdata    (_mmio_io_dma_wdata),
    .io_dma_wstrb    (_mmio_io_dma_wstrb),
    .io_dma_bready        (_mmio_io_dma_bready),
    .io_dma_bvalid        (_soc_io_frontend_bvalid),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_dma_arready       (_soc_io_frontend_arready),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_dma_arvalid       (_mmio_io_dma_arvalid),
    .io_dma_araddr   (_mmio_io_dma_araddr),
    .io_dma_rready        (_mmio_io_dma_rready),
    .io_dma_rvalid        (_soc_io_frontend_rvalid),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_dma_rdata    (_soc_io_frontend_rdata),	// src/main/scala/sim/NutShellSim.scala:28:19
    .io_uart_out_valid     (difftest_uart_out_valid),
    .io_uart_out_ch        (difftest_uart_out_ch),
    .io_uart_in_valid      (difftest_uart_in_valid),
    .io_uart_in_ch         (difftest_uart_in_ch)
  );
  assign difftest_step = 64'h1;	// difftest/src/main/scala/Difftest.scala:395:19, src/main/scala/sim/NutShellSim.scala:26:7
endmodule

